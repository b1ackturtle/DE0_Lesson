module Lesson1(switch, led);
	input switch;
	output led;
	
	assing led=switch;
endmodule
